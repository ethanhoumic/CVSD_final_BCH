// list all paths to your design files
`include "../01_RTL/bch.v"
